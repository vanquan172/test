
                instr_tmp = {seq.RV64A_funct7,seq.RV64A_rs2, seq.RV64A_rs1, seq.RV64A_funct3, seq.RV64A_rd, seq.RV64A_opcode}; 